�P  }@�                                                                                                                                                                 � v�                                ��������������������������������������� v                                  � v                                   ���  c                              ����� �����������������������������������    c                              ��                                  �� �� �                              �����0����������������������������������    �                              ��                                  ������                             _�g���?�����������������������������������  ��                             ���                                 ?��F@���                             ?�?�O����������������������������������?��F@  ��                             ?��F@                                 ?�� ?��@                             �?����������������������������������?��   �@                             ?��    �                             ?���?��@                             �����������������������������������?���  �@                             ?���   �                             �� H���                             {������#���������������������������������� H  ��                             �� H                                  �� (���                             {���������������������������������������� (  ��                             �� (                                       ���                             {��������������������������������������       ��                                                                         ����                             {����� �������������������������������       ��                                                                          ��                               ������ �������������������������������                                                                                    ��                               ������ �������������������������������                                                                                                                      ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                ����������������������                ���������������������������������������                   p                   ����������������������                �@�����������������                �������������������������������������       �          �                   ��@�������������������                ~?� ����������?�������                ~?�������������������������������������� �     �     �|   �                   �W����������?��������                |� ����������������                |�������������������������������������� �   `     ��  �                   ~?� �����������������                x� ��������� p������                x������������������������������������� �   �     ��� �                   |�W���O������ p�����                p� ���_������> �����                p������_������������������������������� D   X     ��� �~                  x������������ ����                `� ����������?0 '�����                `��������������?������������������������ $�  �     �����                  p����S������0 /� ��                @� �� W������� 7�����                @����� W�������������������������������� 7�   V     ����                  `� /��ߩ������� 7��#��                  � ��+������_� �����                  �����+������������������������������?�    +     �� �                  @� ������������ ��c��                  ������������� ���?��                  �����������?�����?�������������������    �    ��  88                    ������������?�������                  ����� J�������������                ;������ J�������������������������������     J�    ? � 0                  8�������?������������                  ������������������                ;�������������������������������������    `    ( �                   8���������������������                  ����� ��������������                ;������ �������������������������������     �    8                     8�������O��������������                  ����� �_�������������                ������ �_������������������������������     �X      	                      ������~���������������                  ����� ���������������                ������ ��������������������������������     �                              �������S��������������                  ����   W��������������                �����   W�������������������������������      V                                ������ߩ��������������                                                        ���������������������������������������                                                                                           �����                                               ���������������                                        �����������    ?��������                          ��                                               ���������������                `                       �����������    ��������                          7�����                                  ���        ���������������                `                       ��������������?��������                 �      o�����                         �        ���        ���������������  �           `                       ����������������������                 i�   <  ������ ��                     h        ���  ��   ���������������  i�   <       ` ��                   ���������������������                 ��   � ������  �                     �        ?���   �   ���������������  ��   �       `  �                   ����������?����� �����                 ``   4�������� ��                     `    4   ?���  ��   ���������������  ``   4�       `  �                   ��������� ?�����������                 �0   pl�� �� ��                     �    p          ��   ���������������  �0   pl          �                   ��������      ��������               ����?��� ������� ��                                    ��   �������������������?���         �                   ���������      ��������               ������� �������?� ���                                 ?� ��� ���������������?�������       ?� ���                 O���������      �� �����               �����?� ���~��������                               ����� ���������������?�����?�       �����                 O���������   �  ��������               ?����������~���?�����                                 ����� ���������������?�������        �����                 ���������  `�  ��������               ?��������������?�����                                 ����� ���������������?�������        �����                 ���������      ��������               8>��p}��������?�����                                  ����� ���������������8>��p}�        �����                 |~��?����      ��������               �،$=�@�������pw����                    �  @       pw���� ����������������،$=�@       pw����                 x>���}��D    ��������                �  @   �����P`7���@                  �  @          `7���@ ��������������� �  @          `7���@                 x?�������    `��w������                                                                               ���������������                                        |��?�������������������                                                                               ���������������                                        ������������������������                                                                               ���������������                                        ������������������������                 a                                       `                     ���������������  a                                     ������������������������                 i�                                      h                     ���������������  i�                                    ������������������������                 ��                                      �                     ���������������  ��                                    ������������������������                 ``                                      `        �           ���������������  ``                                    ������������������������                 �0                                      �        0           ���������������  �0                                    �����������������������               ����      �                                      o�           �������������������                                   ������������������������               ����      �                                      ��          ���������������?����                                   O������������������������               ����      ?�                                    ���          ���������������?����                                   O������������������������               ?����                                           �  �          ���������������?����                                   ����������  ������������               ?����                                           ���          ���������������?����                                  �����������������������               8>��                                            �/�          ���������������8>��                                 |~��?�������������������               ��                                          ���          �����������������                                  x>���������������������                  �                                      �    ���          ���������������   �                                  x?���������������������                                                                �          ���������������                                        |��?������������������                                                                �          ���������������                                        ���������������������                                                                               ���������������                                        ����������������������                                                                               ���������������                                        �����������������������                                                                               ���������������                                        ������������������������                                                                               ���������������                                        ������������������������                                                                               ���������������                                        ������������������������                                                                               ���������������                                        ������������������������                                                                               ���������������                                        ������������������������                                                                               ���������������                                        ������������������������                                                       ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                                      �������������������������                                         �                                      �                                      �           ��                ������ �                                      !                                    � ?  �                                � ?  �      ��                ������H )  �                                � ^� �                                � � �        ��   ��   ��         � � �      ��  �~��        ������� P� �                 ����         � �@ �                                � � ��       ��   ��   ��         � � ��     ��  �~��        ������ `� ��                ����         � �@ ��                               � � ?��  �    ��   ��   ��         � � ?��  �  ��  �~��        ������� P� ?��                ����         � �@ <�  �                            � � |�� �    �?   �    ��         � � |�� �  ��  �~�         ������� � |��                � ��          �@ {~  �                            l m� �~p ��   �?   �    ��         l m� �~p �� ��  �~�         ������l m� �~p                � ��          �@ ��� ��                            a��|8 ��   �    �    ��          a��|8 �� ��  �~�         ������ a��|8                � ��          �@��� ��                           � ���8 ��   �    �    ��         � ���8     ��  �~�         ������� ���8 ��            � ��          �@�{�                                    ��x ��   �    �    ��              ��x     ��  �~�         ������     ��x ��            � ��         � �����                               � ����� 6�h   ��   ��   ��         � ����� 	$� ��  ����        ������� ����� ?��            ����           ��| 	$�                           � ����� ��   ��   ��   ��         � �����     ��  ����        ������� ����� ��            ����           ��                                ���� ��   ��   ��   ��          ����     ��  ����        ������ ���� ��            ����         � ���                               � �����         ?   �    ��         � �����     ��  �~�         ������� �����                � ��         	Y+ �~|                               V ����|         ?   �    ��         V ����|     ��  �~�         ������V ����|                � ��         	�5 ���                               � ����|  �      ?   �    ��         � ����|  �  ��  �~�         ������� ����|                � ��         9Y�+8���  �                            6V������ �    �?   �    �          6V������ �  ��  �~�         ������6V������                � �          I�)5$�x �                            6������ ��   �?   �    �          6������ �� ��  �~�         ������6������                � �          IY)+$��� ��                           6V����� ��   ��   ��   �          6V����� �� ��  �~��        ������6V�����                ���          I�)5$��� ��                           6���� �� ��   ��   ��   �          6���� ��     ��  �~��        ������6���� �� ��            ���          IY)+$ ���                               6V��� ~� ��   ��   ��   �          6V��� ~�     ��  �~��        ������6V��� ~� ��            ���          I�)5$ }��                               6���� ?� -��                           6���� ?� I  ��                ������6���� ?� ?��                           IY)+$ >�� I                            6V��� �� ��                           6V��� ��     ��                ������6V��� �� ��                           I�)5$ �                               7��� �  ��                           7��� �      ��                ������7��� �  ��                           H�)$ �                                7���� �                ��             7���� �      ��    ?���      ������7���� �             ?���             H) $ �                                0 �                    ��             0 �          ��    ?���      ������0 �                 ?���             O�)��                                   0 �                    ��             0 �          ��    ?���      ������0 �                 ?���             H) $                                                           ~�             0 �           ��    ?�~�      ������0 �                 ?�~�             0 �                                                             ~�                         ��    ?�~�      ������0 �                 ?�~�                                                                           ~                             ��    ?�~        ������                     ?�~                                                                               ~                             ��    ?�~        ������                     ?�~                                                                               ~                             ��    ?�~        ������                     ?�~                                                                               ��                           ��     ��      ������                      ��                                                                             ��                           ��     ��      ������                      ��                                                                             ��                           ��     ��      ������                      ��                                                                              �                           ��    �  �      ������                     �  �                                                                              �                           ��    �  �      ������                     �  �                                                                              �                           ��    �  �      ������                     �  �                                                                             ~�                           ��    � ~�      ������                     � ~�                                                                             ~�                           ��    � ~�      ������                     � ~�                                                                             ��                           ��    � ��      ������                     � ��                                                                             ��                           ��    � ��      ������                     � ��                                                                             ��                           ��    � ��      ������                     � ��                                                                                                           ��                ������                                                                                                                                      ��                ������                                                                                                                                      ��                ������                                                                                                   ��   ��                          ��     � ��   ?��������                            ��?��                      �~��� ����?��                         ��   ��                          ��     � ��   ?��������                            ��?��                      �~��� ����?��                         ��   ��                          ��     � ��   ?��������                            ��?��                      �~��� ����?��                         �    ��                          ��     � ��   ?�������                            ��?�                      �~� � ����?�                         �    ��                          ��     � ��   ?�������                            ��?�                      �~� � ����?�                         �    �                           ��     � �    ?�������                            ��?�                      �~� � � ��?�                         �    �                           ��     � �    ?�������                            ��?�                      �~� � � ��?�         �              �    �              ��        ��     � �    ?������� ��                     ��?�                    �~� � � ��?�         @              ��   �             @       ��     � �    ?���������>                    ��?�       ��  �      8p��� � ��?�         @              ��   �              � @    
�   ��     � �    ?�������5�P@*  
�                 ��?�      5�P *          8p��� � ��?�         @              ��   �              �@    �   ��     � �    ?�������?���>  �                 ��?�      ?���>          8p��� � ��?�         �              �    �             1���        ��     � �    ?�������?���                    ��?�      ;�             ?�� � � ��?�         �              �    �             ;� �        ��     � �    ?�������?�@�                    ��?�      ?�@            ?�� � � ��?�      ��    �        �    �              ��6   �   ��     � �    ?������� @�	                    ��?�      �  >  �      ?�� � � ��?�      ?���   �        �    ��             ��6  �   ��     � ��   ?�������?�  I                     ��?�      5��   ?��      �� � ����?�      .���   @        �    ��             ��>  @   ��     � ��   ?�������.�   A                     ��?�      *��  A �@      �� � ����?�      .���   @        ��   ��             ��  @   ��     ����   ?��������.�   A                     ��?��      .��  ] _@@      ���������?��      ��   @        ��   ��             ��  @   ��     ����   ?��������.�   A D@                   ��?��      .��  ] _@@      ���������?��                      ��   ��               �   @   ��     ����   ?��������.��A   @                 ��?��      .�� ]          ���������?��                                              �        ��                ������  �                                    �                                                                           �>        �������������������������  �                                    �  >                                 ?�                                       �>        �������������������������?� �                                   ?��  >                                                                           �       �������������������������
  �                                    �                                                                            ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                                                        ���������������������������������������                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ?� ?� ?� ?� ?� ?� ?������������������@���  ���  ���  ��������������������@   ������     �����������������������@         ������������������������������ ?� ?� ?� ?� ?� ?� ?������������������@���  ���  ���  ��������������������@   ������     �����������������������@         ������������������������������ ?� ?� ?� ?� ?� ?� ?������������������@���  ���  ���  ��������������������@   ������     �����������������������@         ������������������������������ ?� ?� ?� ?� ?� ?� ?������������������@���  ���  ���  ��������������������@   ������     �����������������������@         �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������